module a64dec(input [31:0]i, output v);
    wire [199:0]vtmp;
    assign vtmp[   0] = (i & 32'b00000000000000000000000001110011) == 32'b00000000000000000000000001000011; // esp_0
    assign vtmp[   1] = (i & 32'b00000000000000000000000001011111) == 32'b00000000000000000000000001001111; // esp_1
    assign vtmp[   2] = (i & 32'b00000000000000000000000001011111) == 32'b00000000000000000000000000010111; // esp_2
    assign vtmp[   3] = (i & 32'b00000000000000000010000001111011) == 32'b00000000000000000010000000010011; // esp_3
    assign vtmp[   4] = (i & 32'b00011000000000000000000001001111) == 32'b00001000000000000000000000000111; // esp_4
    assign vtmp[   5] = (i & 32'b00010100000000000000000001001111) == 32'b00000100000000000000000000000111; // esp_5
    assign vtmp[   6] = (i & 32'b00000000000000000010000000111111) == 32'b00000000000000000000000000000011; // esp_6
    assign vtmp[   7] = (i & 32'b00000000000000000110000000111111) == 32'b00000000000000000000000000001111; // esp_7
    assign vtmp[   8] = (i & 32'b00000000000000000111000001001111) == 32'b00000000000000000100000000000111; // esp_8
    assign vtmp[   9] = (i & 32'b00000000000000000010000001111111) == 32'b00000000000000000010000001110011; // esp_9
    assign vtmp[  10] = (i & 32'b00000000000000001111110000000011) == 32'b00000000000000001010000000000010; // esp_10
    assign vtmp[  11] = (i & 32'b00000000000000001111100100000011) == 32'b00000000000000001011100000000010; // esp_11
    assign vtmp[  12] = (i & 32'b00000000000000000111000001110111) == 32'b00000000000000000000000000010011; // esp_12
    assign vtmp[  13] = (i & 32'b00000000000000001111110000100011) == 32'b00000000000000001010110000100010; // esp_13
    assign vtmp[  14] = (i & 32'b00010001111100000000000001001111) == 32'b00000000000000000000000000000111; // esp_14
    assign vtmp[  15] = (i & 32'b11010100000000000011000000101111) == 32'b01000100000000000000000000000111; // esp_15
    assign vtmp[  16] = (i & 32'b10110010000000000100000001101111) == 32'b10000010000000000100000001100011; // esp_16
    assign vtmp[  17] = (i & 32'b11010110000000000111000001011011) == 32'b00000000000000000100000000010011; // esp_17
    assign vtmp[  18] = (i & 32'b10110001110000000100000001101111) == 32'b10000001110000000100000001100011; // esp_18
    assign vtmp[  19] = (i & 32'b11011110000000000111000001010111) == 32'b01000000000000000101000000010011; // esp_19
    assign vtmp[  20] = (i & 32'b10111110000000000111000001010111) == 32'b00000000000000000000000000010011; // esp_20
    assign vtmp[  21] = (i & 32'b11111110000000000100000001110111) == 32'b00000010000000000100000000110011; // esp_21
    assign vtmp[  22] = (i & 32'b11111110000000000011000001110111) == 32'b01100000000000000001000000110011; // esp_22
    assign vtmp[  23] = (i & 32'b11111110000000000101000001110111) == 32'b00100000000000000100000000110011; // esp_23
    assign vtmp[  24] = (i & 32'b11111110000000000011000001110111) == 32'b00100000000000000010000000110011; // esp_24
    assign vtmp[  25] = (i & 32'b11111100000000000110000001111111) == 32'b00001000000000000000000000011011; // esp_25
    assign vtmp[  26] = (i & 32'b11010110000011110110000000101111) == 32'b10010110000000000010000000000111; // esp_26
    assign vtmp[  27] = (i & 32'b11010110000011011110000000101111) == 32'b10010110000000011010000000000111; // esp_27
    assign vtmp[  28] = (i & 32'b11110011111100000100000001101111) == 32'b01100000000000000100000001100011; // esp_28
    assign vtmp[  29] = (i & 32'b11110010000000000100111111101111) == 32'b01100010000000000100000001100011; // esp_29
    assign vtmp[  30] = (i & 32'b11111111110100000100000001101111) == 32'b01100100000100000100000001100011; // esp_30
    assign vtmp[  31] = (i & 32'b11111111110100000100000001101111) == 32'b01101000000100000100000001100011; // esp_31
    assign vtmp[  32] = (i & 32'b00000000000000000110000001011011) == 32'b00000000000000000010000000000011; // esp_32
    assign vtmp[  33] = (i & 32'b00000000000000000101000001011011) == 32'b00000000000000000001000000000011; // esp_33
    assign vtmp[  34] = (i & 32'b00000000000000000001000001101111) == 32'b00000000000000000000000000000011; // esp_34
    assign vtmp[  35] = (i & 32'b00000000000000000100000001011111) == 32'b00000000000000000100000001000011; // esp_35
    assign vtmp[  36] = (i & 32'b00000000000000000100000001011111) == 32'b00000000000000000000000000000011; // esp_36
    assign vtmp[  37] = (i & 32'b00000000000000000111000001011011) == 32'b00000000000000000000000001000011; // esp_37
    assign vtmp[  38] = (i & 32'b00000000000000000011000001101111) == 32'b00000000000000000001000001100011; // esp_38
    assign vtmp[  39] = (i & 32'b00011000000000000100000000111111) == 32'b00000000000000000000000000101111; // esp_39
    assign vtmp[  40] = (i & 32'b11100000000000000000000001101111) == 32'b00000000000000000000000001000011; // esp_40
    assign vtmp[  41] = (i & 32'b11100000000000000111000000101011) == 32'b00000000000000000100000000000011; // esp_41
    assign vtmp[  42] = (i & 32'b11100100000000000010000001101011) == 32'b00000000000000000000000001000011; // esp_42
    assign vtmp[  43] = (i & 32'b11100000000000000101000000101111) == 32'b10100000000000000001000000000111; // esp_43
    assign vtmp[  44] = (i & 32'b01100000000000000111000000101111) == 32'b00000000000000000010000000000111; // esp_44
    assign vtmp[  45] = (i & 32'b10000000000000000111000000111111) == 32'b00000000000000000111000000010111; // esp_45
    assign vtmp[  46] = (i & 32'b01000000000000000111000000111111) == 32'b01000000000000000111000000010111; // esp_46
    assign vtmp[  47] = (i & 32'b11000100000000000001000000111111) == 32'b10000100000000000000000000010111; // esp_47
    assign vtmp[  48] = (i & 32'b10100000000000000011000000111111) == 32'b10000000000000000010000000010111; // esp_48
    assign vtmp[  49] = (i & 32'b11111000000000000010000001101011) == 32'b10100000000000000000000001000011; // esp_49
    assign vtmp[  50] = (i & 32'b11110000000000000110000001101011) == 32'b00010000000000000000000001000011; // esp_50
    assign vtmp[  51] = (i & 32'b10111100000000000100000001101011) == 32'b00101000000000000000000000000011; // esp_51
    assign vtmp[  52] = (i & 32'b11111100000000000000000001011011) == 32'b00000000000000000000000000010011; // esp_52
    assign vtmp[  53] = (i & 32'b11011000000000000100000001110111) == 32'b00001000000000000000000000100111; // esp_53
    assign vtmp[  54] = (i & 32'b10110000000000000110000000111111) == 32'b00000000000000000010000000101111; // esp_54
    assign vtmp[  55] = (i & 32'b11111100000000000000000000101111) == 32'b00100100000000000000000000000111; // esp_55
    assign vtmp[  56] = (i & 32'b11001100000000000110000000101111) == 32'b10000100000000000010000000000111; // esp_56
    assign vtmp[  57] = (i & 32'b11110100000000000010000000101111) == 32'b01100100000000000000000000000111; // esp_57
    assign vtmp[  58] = (i & 32'b01101000000000000111000000101111) == 32'b00101000000000000011000000000111; // esp_58
    assign vtmp[  59] = (i & 32'b11111000000000000001000000101111) == 32'b00101000000000000000000000000111; // esp_59
    assign vtmp[  60] = (i & 32'b01011100000000000011000000101111) == 32'b00001000000000000000000000000111; // esp_60
    assign vtmp[  61] = (i & 32'b11100000000000000111000000101111) == 32'b01100000000000000100000000000111; // esp_61
    assign vtmp[  62] = (i & 32'b11000100000000000110000000111111) == 32'b11000000000000000110000000010111; // esp_62
    assign vtmp[  63] = (i & 32'b10110000000000000011000000111111) == 32'b10110000000000000001000000010111; // esp_63
    assign vtmp[  64] = (i & 32'b10001100000000000011000000111111) == 32'b10000000000000000001000000010111; // esp_64
    assign vtmp[  65] = (i & 32'b10001100000000000011000000111111) == 32'b10001100000000000010000000010111; // esp_65
    assign vtmp[  66] = (i & 32'b00010000111100000000000000111111) == 32'b00000000000000000000000000000111; // esp_66
    assign vtmp[  67] = (i & 32'b00110010000000000111000001001111) == 32'b00100010000000000000000000000011; // esp_67
    assign vtmp[  68] = (i & 32'b01111000000000000101000000101111) == 32'b00100000000000000000000000000011; // esp_68
    assign vtmp[  69] = (i & 32'b11011000000000000100000001101111) == 32'b00001000000000000000000001000011; // esp_69
    assign vtmp[  70] = (i & 32'b11011100000000000110000001101011) == 32'b00000100000000000000000001000011; // esp_70
    assign vtmp[  71] = (i & 32'b11010100000000000111000001101011) == 32'b00000000000000000001000001000011; // esp_71
    assign vtmp[  72] = (i & 32'b10111110000000000100000001011011) == 32'b00000000000000000100000000010011; // esp_72
    assign vtmp[  73] = (i & 32'b11111100000000000000000001111011) == 32'b01001000000000000000000000010011; // esp_73
    assign vtmp[  74] = (i & 32'b11101000000000000110000000111111) == 32'b00001000000000000010000000101111; // esp_74
    assign vtmp[  75] = (i & 32'b10111100000000000110000000101111) == 32'b10010100000000000010000000000111; // esp_75
    assign vtmp[  76] = (i & 32'b11110010000000000110000000101111) == 32'b01110010000000000010000000000111; // esp_76
    assign vtmp[  77] = (i & 32'b11001010000000000111000000101111) == 32'b01000000000000000011000000000111; // esp_77
    assign vtmp[  78] = (i & 32'b11111000000000000100000000111111) == 32'b00111000000000000100000000010111; // esp_78
    assign vtmp[  79] = (i & 32'b01111100000000000100000000111111) == 32'b00000000000000000000000000010111; // esp_79
    assign vtmp[  80] = (i & 32'b11011000000000000110000000111111) == 32'b10000000000000000100000000010111; // esp_80
    assign vtmp[  81] = (i & 32'b11100100000000000110000000111111) == 32'b01100100000000000100000000010111; // esp_81
    assign vtmp[  82] = (i & 32'b11101100000000000001000000111111) == 32'b01100000000000000001000000010111; // esp_82
    assign vtmp[  83] = (i & 32'b11011000000000000011000000111111) == 32'b01010000000000000011000000010111; // esp_83
    assign vtmp[  84] = (i & 32'b11001100000000000011000000111111) == 32'b01000100000000000011000000010111; // esp_84
    assign vtmp[  85] = (i & 32'b10110100000000000011000000111111) == 32'b00110000000000000011000000010111; // esp_85
    assign vtmp[  86] = (i & 32'b10101100000000000011000000111111) == 32'b10101100000000000001000000010111; // esp_86
    assign vtmp[  87] = (i & 32'b11100100000000000011000000111111) == 32'b11000000000000000001000000010111; // esp_87
    assign vtmp[  88] = (i & 32'b01110100000000000011000000111111) == 32'b00100000000000000001000000010111; // esp_88
    assign vtmp[  89] = (i & 32'b11101000000000000011000000111111) == 32'b00100000000000000010000000010111; // esp_89
    assign vtmp[  90] = (i & 32'b11011000000000000011000000111111) == 32'b11010000000000000010000000010111; // esp_90
    assign vtmp[  91] = (i & 32'b11010100000000000011000000111111) == 32'b11000000000000000010000000010111; // esp_91
    assign vtmp[  92] = (i & 32'b11011000000000000011000000111111) == 32'b01010000000000000000000000010111; // esp_92
    assign vtmp[  93] = (i & 32'b00111100000000000011000000111111) == 32'b00010100000000000000000000010111; // esp_93
    assign vtmp[  94] = (i & 32'b01110100000000000011000000111111) == 32'b00110000000000000000000000010111; // esp_94
    assign vtmp[  95] = (i & 32'b11010010000000000011000000111111) == 32'b01000000000000000000000000010111; // esp_95
    assign vtmp[  96] = (i & 32'b11100010000000000111000001001111) == 32'b00100010000000000000000000000011; // esp_96
    assign vtmp[  97] = (i & 32'b00111010000000000111000001001111) == 32'b00110000000000000000000000000011; // esp_97
    assign vtmp[  98] = (i & 32'b11110110000000000010000000011111) == 32'b00000010000000000010000000010011; // esp_98
    assign vtmp[  99] = (i & 32'b10111110000000000111000001001011) == 32'b00101000000000000001000000000011; // esp_99
    assign vtmp[ 100] = (i & 32'b11111100000000000101000001101011) == 32'b00001100000000000001000001000011; // esp_100
    assign vtmp[ 101] = (i & 32'b11110110000000000100000001111011) == 32'b00000010000000000100000000110011; // esp_101
    assign vtmp[ 102] = (i & 32'b11111000000000000011000000111111) == 32'b00101000000000000000000000101111; // esp_102
    assign vtmp[ 103] = (i & 32'b11010110000000000111000000101111) == 32'b01010100000000000011000000000111; // esp_103
    assign vtmp[ 104] = (i & 32'b11011100000000000111000000101111) == 32'b11001100000000000001000000000111; // esp_104
    assign vtmp[ 105] = (i & 32'b00111110000000000111000000101111) == 32'b00011110000000000010000000000111; // esp_105
    assign vtmp[ 106] = (i & 32'b11111110000000000000000000111111) == 32'b10000000000000000000000000010111; // esp_106
    assign vtmp[ 107] = (i & 32'b11011100000000000110000000111111) == 32'b10011100000000000100000000010111; // esp_107
    assign vtmp[ 108] = (i & 32'b11111000000000000110000000111111) == 32'b11000000000000000000000000010111; // esp_108
    assign vtmp[ 109] = (i & 32'b11110010000000000101000000111111) == 32'b01100010000000000000000000010111; // esp_109
    assign vtmp[ 110] = (i & 32'b10110110000000000011000000111111) == 32'b00010100000000000000000000010111; // esp_110
    assign vtmp[ 111] = (i & 32'b11111000000000000111000001001111) == 32'b01010000000000000000000000000011; // esp_111
    assign vtmp[ 112] = (i & 32'b11110100000000000111000001001111) == 32'b01010100000000000000000000000011; // esp_112
    assign vtmp[ 113] = (i & 32'b11101010000000000111000000101111) == 32'b10100010000000000000000000000011; // esp_113
    assign vtmp[ 114] = (i & 32'b11101001110000000000000001101111) == 32'b11000000000000000000000001000011; // esp_114
    assign vtmp[ 115] = (i & 32'b11011100000000000110000001101111) == 32'b01000000000000000100000000000011; // esp_115
    assign vtmp[ 116] = (i & 32'b11110100000000000111000000011111) == 32'b00000000000000000111000000010011; // esp_116
    assign vtmp[ 117] = (i & 32'b11110110000000000001000000111111) == 32'b00000010000000000001000000110011; // esp_117
    assign vtmp[ 118] = (i & 32'b11111110000000000011000001011011) == 32'b01001000000000000001000000010011; // esp_118
    assign vtmp[ 119] = (i & 32'b11111010000000000111000000011111) == 32'b10000010000000000010000000010111; // esp_119
    assign vtmp[ 120] = (i & 32'b11110010000000000111000000111111) == 32'b10110010000000000010000000110111; // esp_120
    assign vtmp[ 121] = (i & 32'b11101010000000000111000000111111) == 32'b10101010000000000010000000110111; // esp_121
    assign vtmp[ 122] = (i & 32'b11011110000000000110000000111111) == 32'b01011100000000000100000000010111; // esp_122
    assign vtmp[ 123] = (i & 32'b11010011011100000000000000111111) == 32'b00000010000000000000000000000111; // esp_123
    assign vtmp[ 124] = (i & 32'b01110011011100000000000000111111) == 32'b01100010000000000000000000000111; // esp_124
    assign vtmp[ 125] = (i & 32'b11111110000000000011000001010111) == 32'b00000000000000000001000000010011; // esp_125
    assign vtmp[ 126] = (i & 32'b11011110000000000111000001001111) == 32'b01011110000000000000000000000011; // esp_126
    assign vtmp[ 127] = (i & 32'b10111001111000000000000001101111) == 32'b00000000010000000000000001000011; // esp_127
    assign vtmp[ 128] = (i & 32'b11110110000000000111000000011111) == 32'b00100000000000000010000000010011; // esp_128
    assign vtmp[ 129] = (i & 32'b11111010000000000101000000111111) == 32'b00001010000000000101000000110011; // esp_129
    assign vtmp[ 130] = (i & 32'b11101111100000000100000001111011) == 32'b00000000000000000000000000010011; // esp_130
    assign vtmp[ 131] = (i & 32'b01111100000011000111000000101111) == 32'b01001000000001000001000000000111; // esp_131
    assign vtmp[ 132] = (i & 32'b01111100000011000111000000101111) == 32'b01001000000010000001000000000111; // esp_132
    assign vtmp[ 133] = (i & 32'b01111100000001100111000000101111) == 32'b01001000000000000001000000000111; // esp_133
    assign vtmp[ 134] = (i & 32'b01111100000001010111000000101111) == 32'b01001000000000010001000000000111; // esp_134
    assign vtmp[ 135] = (i & 32'b00111100000011100111000000101111) == 32'b00001000000000100010000000000111; // esp_135
    assign vtmp[ 136] = (i & 32'b00111100000011010111000000101111) == 32'b00001000000000010010000000000111; // esp_136
    assign vtmp[ 137] = (i & 32'b00111100000011010111000000101111) == 32'b00001000000001000010000000000111; // esp_137
    assign vtmp[ 138] = (i & 32'b00111100000010011111000000101111) == 32'b00001000000000010010000000000111; // esp_138
    assign vtmp[ 139] = (i & 32'b11011110000000000111000000111111) == 32'b10001010000000000010000000110111; // esp_139
    assign vtmp[ 140] = (i & 32'b11111110000000000011000001110111) == 32'b00000010000000000000000000110011; // esp_140
    assign vtmp[ 141] = (i & 32'b01111101111000000000000001101111) == 32'b01000000001000000000000001000011; // esp_141
    assign vtmp[ 142] = (i & 32'b01111101111000000000000001101111) == 32'b01000100000000000000000001000011; // esp_142
    assign vtmp[ 143] = (i & 32'b01111011110100000000000001101111) == 32'b01000000000100000000000001000011; // esp_143
    assign vtmp[ 144] = (i & 32'b01111011110100000000000001101111) == 32'b01000010000000000000000001000011; // esp_144
    assign vtmp[ 145] = (i & 32'b10111001111100000000000001101111) == 32'b00011000000000000000000001000011; // esp_145
    assign vtmp[ 146] = (i & 32'b11111111000000000100000001101111) == 32'b00110001000000000000000000000011; // esp_146
    assign vtmp[ 147] = (i & 32'b11101111011000000100000001111011) == 32'b00000000000000000000000000010011; // esp_147
    assign vtmp[ 148] = (i & 32'b01111011011100000110000001010111) == 32'b01100010000000000000000000000111; // esp_148
    assign vtmp[ 149] = (i & 32'b11100001111100000110000000111111) == 32'b00000000000000000010000000101111; // esp_149
    assign vtmp[ 150] = (i & 32'b01011100000001111111000000101111) == 32'b01001100000000000001000000000111; // esp_150
    assign vtmp[ 151] = (i & 32'b00111100000011110111000000101111) == 32'b00000000000010000010000000000111; // esp_151
    assign vtmp[ 152] = (i & 32'b11111110000000000011000001111111) == 32'b00001000000000000000000000111011; // esp_152
    assign vtmp[ 153] = (i & 32'b10111111101100000000000001101111) == 32'b00000000001000000000000001000011; // esp_153
    assign vtmp[ 154] = (i & 32'b10111111011100000000000001101111) == 32'b00000100000000000000000001000011; // esp_154
    assign vtmp[ 155] = (i & 32'b11011111011100000111000001001011) == 32'b00000010000000000000000000000011; // esp_155
    assign vtmp[ 156] = (i & 32'b10111111111100000000000001111011) == 32'b00101000011100000000000000010011; // esp_156
    assign vtmp[ 157] = (i & 32'b11110011111100000011000001001111) == 32'b00000010101100000000000000000111; // esp_157
    assign vtmp[ 158] = (i & 32'b10111100000011110111000000101111) == 32'b00001100000000100001000000000111; // esp_158
    assign vtmp[ 159] = (i & 32'b01111100000001111111000000101111) == 32'b01001000000001101001000000000111; // esp_159
    assign vtmp[ 160] = (i & 32'b00111110000001111111000000101111) == 32'b00000010000000000010000000000111; // esp_160
    assign vtmp[ 161] = (i & 32'b11011010000011100111000000111111) == 32'b10000010000000000010000000110111; // esp_161
    assign vtmp[ 162] = (i & 32'b11010110000001110111000000111111) == 32'b10000010000000000010000000110111; // esp_162
    assign vtmp[ 163] = (i & 32'b10111100000011110101000000111111) == 32'b00010000000000010000000000010111; // esp_163
    assign vtmp[ 164] = (i & 32'b10111100000011101101000000111111) == 32'b00010000000000001000000000010111; // esp_164
    assign vtmp[ 165] = (i & 32'b10110101111100000011000000111111) == 32'b00010100000000000000000000010111; // esp_165
    assign vtmp[ 166] = (i & 32'b11011001111100000111000001001111) == 32'b11000000000000000001000001000011; // esp_166
    assign vtmp[ 167] = (i & 32'b11110111111000000100000001101111) == 32'b01100000000000000100000001100011; // esp_167
    assign vtmp[ 168] = (i & 32'b11011011111000000111000000101111) == 32'b11010000000000000000000000000011; // esp_168
    assign vtmp[ 169] = (i & 32'b11001011111100000111000000101111) == 32'b11000010000100000000000000000011; // esp_169
    assign vtmp[ 170] = (i & 32'b11001101111100000111000000101111) == 32'b11000000000000000000000000000011; // esp_170
    assign vtmp[ 171] = (i & 32'b11001011111100000111000000101111) == 32'b11000000000000000000000000000011; // esp_171
    assign vtmp[ 172] = (i & 32'b11111111101000000010000001101111) == 32'b01100000000000000000000000000011; // esp_172
    assign vtmp[ 173] = (i & 32'b11010101111100000110000001101111) == 32'b01000001100000000100000000000011; // esp_173
    assign vtmp[ 174] = (i & 32'b11110111111100000000000000111111) == 32'b00000000111100000000000000010011; // esp_174
    assign vtmp[ 175] = (i & 32'b01111111111100000110000000111011) == 32'b01000010000000000110000000010011; // esp_175
    assign vtmp[ 176] = (i & 32'b10111111111100000101000000111011) == 32'b00000010000000000101000000010011; // esp_176
    assign vtmp[ 177] = (i & 32'b11011111111100000110000000101111) == 32'b01011110000000000010000000000111; // esp_177
    assign vtmp[ 178] = (i & 32'b01110110000011111111000000101111) == 32'b01000010000000000001000000000111; // esp_178
    assign vtmp[ 179] = (i & 32'b11011010000001111111000000111111) == 32'b10000010000000000010000000110111; // esp_179
    assign vtmp[ 180] = (i & 32'b11011101111100000110000000111111) == 32'b01011100000000000100000000010111; // esp_180
    assign vtmp[ 181] = (i & 32'b10111100000011111101000000111111) == 32'b00010000000010000000000000010111; // esp_181
    assign vtmp[ 182] = (i & 32'b11011111111100000100000001101111) == 32'b00010000000000000000000000000011; // esp_182
    assign vtmp[ 183] = (i & 32'b11111010000000000100111111011111) == 32'b00010010000000000000000001010011; // esp_183
    assign vtmp[ 184] = (i & 32'b10111010000000000100111111111111) == 32'b00100010000000000000000001110011; // esp_184
    assign vtmp[ 185] = (i & 32'b11011110000011011111000001111011) == 32'b10000110000000011010000001110011; // esp_185
    assign vtmp[ 186] = (i & 32'b11111111111000000110000001110111) == 32'b01100000000000000000000000010011; // esp_186
    assign vtmp[ 187] = (i & 32'b11111111110100000110000001110111) == 32'b01100000000000000000000000010011; // esp_187
    assign vtmp[ 188] = (i & 32'b11111111011100000111000001001111) == 32'b11000010000000000001000001000011; // esp_188
    assign vtmp[ 189] = (i & 32'b10111101111101111101000000111111) == 32'b00010000000000001000000000010111; // esp_189
    assign vtmp[ 190] = (i & 32'b11111111111000000111111110110111) == 32'b00000000000000000010000000000111; // esp_190
    assign vtmp[ 191] = (i & 32'b11111111110100000111111110110111) == 32'b00000000000000000010000000000111; // esp_191
    assign vtmp[ 192] = (i & 32'b11111111101100000111111110110111) == 32'b00000000000000000010000000000111; // esp_192
    assign vtmp[ 193] = (i & 32'b11111111111011111100111110011111) == 32'b00000000000000000000000000010011; // esp_193
    assign vtmp[ 194] = (i & 32'b11111110111111111100111110011111) == 32'b00000000110100000000000000010011; // esp_194
    assign vtmp[ 195] = (i & 32'b11111101111011111100111111011111) == 32'b00010000010000000000000001010011; // esp_195
    assign vtmp[ 196] = (i & 32'b11111111111011111100111111011111) == 32'b00011000000000000000000001010011; // esp_196
    assign vtmp[ 197] = (i & 32'b11011111111111111100111111111111) == 32'b00010000001000000000000001110011; // esp_197
    assign vtmp[ 198] = (i & 32'b10111111111111111100111111111111) == 32'b00110000001000000000000001110011; // esp_198
    assign vtmp[ 199] = (i & 32'b11111111111111111100111111111111) == 32'b01111011001000000000000001110011; // esp_199
    assign v = |vtmp;
endmodule
